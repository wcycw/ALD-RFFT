
`timescale 1ns/1ps
`define HALF_CLOCK_PERIOD #1

module Testbench();

parameter WIDTH = 16;
reg	[WIDTH - 1 : 0] ram [0 : 256];
reg [WIDTH - 1 : 0] Dout0, Dout1, Dout2, Dout3;
reg [WIDTH - 1 : 0] Din0, Din1, Din2, Din3;
reg [5 : 0] addr_I;
reg clk, reset_n;
reg Einput, Ewrite;
reg done;

rfft rfft0(.Clk(clk), .Reset_n(reset_n), .done(done), .Din0(Din0), .Din1(Din1), .Din2(Din2), .Din3(Din3), .Dout0(Dout0), .Dout1(Dout1), .Dout2(Dout2), .Dout3(Dout3), .Addr(addr_I), .Input(Einput), .Write(Ewrite));

always begin
	`HALF_CLOCK_PERIOD;
	clk = ~clk;
end

initial begin

clk = 0;
resetn = 0;
ram[0] = {8'd1,8'b00000000};
ram[1] = {8'd1,8'b00000000};
ram[2] = {8'd4,8'b00000000};
ram[3] = {8'd1,8'b00000000};
ram[4] = {8'd1,8'b00000000};
ram[5] = {8'd7,8'b00000000};
ram[6] = {8'd1,8'b00000000};
ram[7] = {8'd1,8'b00000000};
ram[8] = {8'd2,8'b00000000};
ram[9] = {8'd5,8'b00000000};
ram[10] = {8'd6,8'b00000000};
ram[11] = {8'd5,8'b00000000};
ram[12] = {8'd1,8'b00000000};
ram[13] = {8'd1,8'b00000000};
ram[14] = {8'd1,8'b00000000};
ram[15] = {8'd1,8'b00000000};
ram[16] = {8'd1,8'b00000000};
ram[17] = {8'd1,8'b00000000};
ram[18] = {8'd2,8'b00000000};
ram[19] = {8'd9,8'b00000000};
ram[20] = {8'd7,8'b00000000};
ram[21] = {8'd8,8'b00000000};
ram[22] = {8'd1,8'b00000000};
ram[23] = {8'd5,8'b00000000};
ram[24] = {8'd3,8'b00000000};
ram[25] = {8'd1,8'b00000000};
ram[26] = {8'd9,8'b00000000};
ram[27] = {8'd5,8'b00000000};
ram[28] = {8'd1,8'b00000000};
ram[29] = {8'd9,8'b00000000};
ram[30] = {8'd1,8'b00000000};
ram[31] = {8'd1,8'b00000000};
ram[32] = {8'd1,8'b00000000};
ram[33] = {8'd3,8'b00000000};
ram[34] = {8'd6,8'b00000000};
ram[35] = {8'd5,8'b00000000};
ram[36] = {8'd4,8'b00000000};
ram[37] = {8'd1,8'b00000000};
ram[38] = {8'd1,8'b00000000};
ram[39] = {8'd2,8'b00000000};
ram[40] = {8'd2,8'b00000000};
ram[41] = {8'd8,8'b00000000};
ram[42] = {8'd8,8'b00000000};
ram[43] = {8'd1,8'b00000000};
ram[44] = {8'd2,8'b00000000};
ram[45] = {8'd1,8'b00000000};
ram[46] = {8'd4,8'b00000000};
ram[47] = {8'd1,8'b00000000};
ram[48] = {8'd3,8'b00000000};
ram[49] = {8'd9,8'b00000000};
ram[50] = {8'd1,8'b00000000};
ram[51] = {8'd7,8'b00000000};
ram[52] = {8'd1,8'b00000000};
ram[53] = {8'd2,8'b00000000};
ram[54] = {8'd5,8'b00000000};
ram[55] = {8'd7,8'b00000000};
ram[56] = {8'd6,8'b00000000};
ram[57] = {8'd2,8'b00000000};
ram[58] = {8'd5,8'b00000000};
ram[59] = {8'd8,8'b00000000};
ram[60] = {8'd3,8'b00000000};
ram[61] = {8'd2,8'b00000000};
ram[62] = {8'd3,8'b00000000};
ram[63] = {8'd1,8'b00000000};
ram[64] = {8'd7,8'b00000000};
ram[65] = {8'd4,8'b00000000};
ram[66] = {8'd2,8'b00000000};
ram[67] = {8'd1,8'b00000000};
ram[68] = {8'd8,8'b00000000};
ram[69] = {8'd6,8'b00000000};
ram[70] = {8'd1,8'b00000000};
ram[71] = {8'd3,8'b00000000};
ram[72] = {8'd4,8'b00000000};
ram[73] = {8'd4,8'b00000000};
ram[74] = {8'd4,8'b00000000};
ram[75] = {8'd5,8'b00000000};
ram[76] = {8'd2,8'b00000000};
ram[77] = {8'd3,8'b00000000};
ram[78] = {8'd9,8'b00000000};
ram[79] = {8'd1,8'b00000000};
ram[80] = {8'd1,8'b00000000};
ram[81] = {8'd3,8'b00000000};
ram[82] = {8'd1,8'b00000000};
ram[83] = {8'd1,8'b00000000};
ram[84] = {8'd8,8'b00000000};
ram[85] = {8'd4,8'b00000000};
ram[86] = {8'd3,8'b00000000};
ram[87] = {8'd5,8'b00000000};
ram[88] = {8'd5,8'b00000000};
ram[89] = {8'd2,8'b00000000};
ram[90] = {8'd1,8'b00000000};
ram[91] = {8'd5,8'b00000000};
ram[92] = {8'd2,8'b00000000};
ram[93] = {8'd3,8'b00000000};
ram[94] = {8'd3,8'b00000000};
ram[95] = {8'd1,8'b00000000};
ram[96] = {8'd4,8'b00000000};
ram[97] = {8'd2,8'b00000000};
ram[98] = {8'd1,8'b00000000};
ram[99] = {8'd7,8'b00000000};
ram[100] = {8'd2,8'b00000000};
ram[101] = {8'd6,8'b00000000};
ram[102] = {8'd2,8'b00000000};
ram[103] = {8'd2,8'b00000000};
ram[104] = {8'd2,8'b00000000};
ram[105] = {8'd2,8'b00000000};
ram[106] = {8'd9,8'b00000000};
ram[107] = {8'd5,8'b00000000};
ram[108] = {8'd5,8'b00000000};
ram[109] = {8'd2,8'b00000000};
ram[110] = {8'd6,8'b00000000};
ram[111] = {8'd3,8'b00000000};
ram[112] = {8'd4,8'b00000000};
ram[113] = {8'd7,8'b00000000};
ram[114] = {8'd5,8'b00000000};
ram[115] = {8'd5,8'b00000000};
ram[116] = {8'd7,8'b00000000};
ram[117] = {8'd6,8'b00000000};
ram[118] = {8'd6,8'b00000000};
ram[119] = {8'd7,8'b00000000};
ram[120] = {8'd9,8'b00000000};
ram[121] = {8'd7,8'b00000000};
ram[122] = {8'd3,8'b00000000};
ram[123] = {8'd7,8'b00000000};
ram[124] = {8'd2,8'b00000000};
ram[125] = {8'd6,8'b00000000};
ram[126] = {8'd6,8'b00000000};
ram[127] = {8'd3,8'b00000000};
ram[128] = {8'd3,8'b00000000};
ram[129] = {8'd4,8'b00000000};
ram[130] = {8'd7,8'b00000000};
ram[131] = {8'd5,8'b00000000};
ram[132] = {8'd8,8'b00000000};
ram[133] = {8'd9,8'b00000000};
ram[134] = {8'd9,8'b00000000};
ram[135] = {8'd4,8'b00000000};
ram[136] = {8'd1,8'b00000000};
ram[137] = {8'd8,8'b00000000};
ram[138] = {8'd2,8'b00000000};
ram[139] = {8'd1,8'b00000000};
ram[140] = {8'd1,8'b00000000};
ram[141] = {8'd2,8'b00000000};
ram[142] = {8'd2,8'b00000000};
ram[143] = {8'd8,8'b00000000};
ram[144] = {8'd7,8'b00000000};
ram[145] = {8'd1,8'b00000000};
ram[146] = {8'd1,8'b00000000};
ram[147] = {8'd1,8'b00000000};
ram[148] = {8'd1,8'b00000000};
ram[149] = {8'd1,8'b00000000};
ram[150] = {8‘d14,8'b00000000};
ram[151] = {8'd1,8'b00000000};
ram[152] = {8'd2,8'b00000000};
ram[153] = {8'd2,8'b00000000};
ram[154] = {8'd1,8'b00000000};
ram[155] = {8'd4,8'b00000000};
ram[156] = {8'd13,8'b00000000};
ram[157] = {8'd2,8'b00000000};
ram[158] = {8'd1,8'b00000000};
ram[159] = {8'd5,8'b00000000};
ram[160] = {8'd3,8'b00000000};
ram[161] = {8'd5,8'b00000000};
ram[162] = {8'd2,8'b00000000};
ram[163] = {8'd1,8'b00000000};
ram[164] = {8'd1,8'b00000000};
ram[165] = {8'd8,8'b00000000};
ram[166] = {8'd7,8'b00000000};
ram[167] = {8'd3,8'b00000000};
ram[168] = {8'd8,8'b00000000};
ram[169] = {8'd5,8'b00000000};
ram[170] = {8'd1,8'b00000000};
ram[171] = {8'd8,8'b00000000};
ram[172] = {8'd3,8'b00000000};
ram[173] = {8'd1,8'b00000000};
ram[174] = {8'd1,8'b00000000};
ram[175] = {8'd7,8'b00000000};
ram[176] = {8'd1,8'b00000000};
ram[177] = {8'd2,8'b00000000};
ram[178] = {8'd2,8'b00000000};
ram[179] = {8'd1,8'b00000000};
ram[180] = {8'd1,8'b00000000};
ram[181] = {8'd3,8'b00000000};
ram[182] = {8'd2,8'b00000000};
ram[183] = {8'd9,8'b00000000};
ram[184] = {8'd1,8'b00000000};
ram[185] = {8'd2,8'b00000000};
ram[186] = {8'd1,8'b00000000};
ram[187] = {8'd2,8'b00000000};
ram[188] = {8'd1,8'b00000000};
ram[189] = {8'd6,8'b00000000};
ram[190] = {8'd8,8'b00000000};
ram[191] = {8'd1,8'b00000000};
ram[192] = {8'd3,8'b00000000};
ram[193] = {8'd1,8'b00000000};
ram[194] = {8'd1,8'b00000000};
ram[195] = {8'd1,8'b00000000};
ram[196] = {8'd9,8'b00000000};
ram[197] = {8'd0,8'b00000000};
ram[198] = {8'd4,8'b00000000};
ram[199] = {8'd1,8'b00000000};
ram[200] = {8'd1,8'b00000000};
ram[201] = {8'd2,8'b00000000};
ram[202] = {8'd2,8'b00000000};
ram[203] = {8'd1,8'b00000000};
ram[204] = {8'd1,8'b00000000};
ram[205] = {8'd3,8'b00000000};
ram[206] = {8'd8,8'b00000000};
ram[207] = {8'd1,8'b00000000};
ram[208] = {8'd1,8'b00000000};
ram[209] = {8'd6,8'b00000000};
ram[210] = {8'd3,8'b00000000};
ram[211] = {8'd2,8'b00000000};
ram[212] = {8'd8,8'b00000000};
ram[213] = {8'd1,8'b00000000};
ram[214] = {8'd1,8'b00000000};
ram[215] = {8'd1,8'b00000000};
ram[216] = {8'd1,8'b00000000};
ram[217] = {8'd7,8'b00000000};
ram[218] = {8'd1,8'b00000000};
ram[219] = {8'd5,8'b00000000};
ram[220] = {8'd1,8'b00000000};
ram[221] = {8'd1,8'b00000000};
ram[222] = {8'd1,8'b00000000};
ram[223] = {8'd8,8'b00000000};
ram[224] = {8'd3,8'b00000000};
ram[225] = {8'd2,8'b00000000};
ram[226] = {8'd4,8'b00000000};
ram[227] = {8'd2,8'b00000000};
ram[228] = {8'd1,8'b00000000};
ram[229] = {8'd2,8'b00000000};
ram[230] = {8'd3,8'b00000000};
ram[231] = {8'd9,8'b00000000};
ram[232] = {8'd1,8'b00000000};
ram[233] = {8'd1,8'b00000000};
ram[234] = {8'd8,8'b00000000};
ram[235] = {8'd9,8'b00000000};
ram[236] = {8'd1,8'b00000000};
ram[237] = {8'd1,8'b00000000};
ram[238] = {8'd3,8'b00000000};
ram[239] = {8'd3,8'b00000000};
ram[240] = {8'd9,8'b00000000};
ram[241] = {8'd1,8'b00000000};
ram[242] = {8'd8,8'b00000000};
ram[243] = {8'd1,8'b00000000};
ram[244] = {8'd1,8'b00000000};
ram[245] = {8'd1,8'b00000000};
ram[246] = {8'd6,8'b00000000};
ram[247] = {8'd1,8'b00000000};
ram[248] = {8'd2,8'b00000000};
ram[249] = {8'd1,8'b00000000};
ram[250] = {8'd7,8'b00000000};
ram[251] = {8'd7,8'b00000000};
ram[252] = {8'd8,8'b00000000};
ram[253] = {8'd1,8'b00000000};
ram[254] = {8'd6,8'b00000000};
ram[255] = {8'd6,8'b00000000};
@(posedge clk);

@(negedge clk);
reset_n = 1;

@(posedge clk);
Einput = 1;
Eoutput = 0;
for (i=0 ; i<64 ; i=i+1)
begin
	addr_I= i;
	Din0 = ram[i*4];
	Din1 = ram[i*4 + 1];
	Din2 = ram[i*4 + 2];
	Din3 = ram[i*4 + 3];
	@(posedge clk);
end

Einput = 0;

@(posedge done);
@(posedge clk);
Ewrite = 0;

for (i=0 ; i<64 ; i=i+1)
begin
	addr_I= i;
	ram[i*4] = Dout0 ;
	ram[i*4 + 1] = Dout1 ;
	ram[i*4 + 2] = Dout2 ;
	ram[i*4 + 3] = Dout3 ;
	@(posedge clk);
end



end
