`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:37:05 03/10/2017 
// Design Name: 
// Module Name:    bram_dual 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bram_duel_T(
	Clk, En, We_A, Addr_A,  DI_A,  DO_A, We_B, Addr_B,  DI_B,  DO_B
    );
parameter WIDTH = 32;

input 		Clk;
input 		En;
input 		We_A;
input		We_B;
input 		[7 : 0]		Addr_A;

input 		[2 * WIDTH - 1 : 0]	DI_A;
output 		[2 * WIDTH - 1 : 0]	DO_A;
reg	 	[2 * WIDTH - 1 : 0]	DO_A;

input 		[7 : 0]		Addr_B;

input 		[2 * WIDTH - 1 : 0]	DI_B;
output 		[2 * WIDTH - 1 : 0]	DO_B;
reg	 	[2 * WIDTH - 1 : 0]	DO_B;

reg 		[2 * WIDTH - 1 : 0]	ram 	 [0 : 255];

initial begin
ram[ 0 ]= 64'b 0000000000000001000000000000000000000000000000000000000000000000;
ram[ 1 ]= 64'b 0000000000000000111111111110110000000000000000000000011001001000;
ram[ 2 ]= 64'b 0000000000000000111111111011000100000000000000000000110010001111;
ram[ 3 ]= 64'b 0000000000000000111111110100111000000000000000000001001011010101;
ram[ 4 ]= 64'b 0000000000000000111111101100010000000000000000000001100100010111;
ram[ 5 ]= 64'b 0000000000000000111111100001001100000000000000000001111101010110;
ram[ 6 ]= 64'b 0000000000000000111111010011101000000000000000000010010110010000;
ram[ 7 ]= 64'b 0000000000000000111111000011101100000000000000000010101111000100;
ram[ 8 ]= 64'b 0000000000000000111110110001010000000000000000000011000111110001;
ram[ 9 ]= 64'b 0000000000000000111110011100011100000000000000000011100000010111;
ram[ 10 ]= 64'b 0000000000000000111110000101001100000000000000000011111000110011;
ram[ 11 ]= 64'b 0000000000000000111101101011101000000000000000000100010001000111;
ram[ 12 ]= 64'b 0000000000000000111101001111101000000000000000000100101001010000;
ram[ 13 ]= 64'b 0000000000000000111100110001010000000000000000000101000001001101;
ram[ 14 ]= 64'b 0000000000000000111100010000100100000000000000000101011000111110;
ram[ 15 ]= 64'b 0000000000000000111011101101100000000000000000000101110000100010;
ram[ 16 ]= 64'b 0000000000000000111011001000001100000000000000000110000111110111;
ram[ 17 ]= 64'b 0000000000000000111010100000100100000000000000000110011110111101;
ram[ 18 ]= 64'b 0000000000000000111001110110101100000000000000000110110101110100;
ram[ 19 ]= 64'b 0000000000000000111001001010101000000000000000000111001100011001;
ram[ 20 ]= 64'b 0000000000000000111000011100010100000000000000000111100010101101;
ram[ 21 ]= 64'b 0000000000000000110111101011111000000000000000000111111000101110;
ram[ 22 ]= 64'b 0000000000000000110110111001010000000000000000001000001110011100;
ram[ 23 ]= 64'b 0000000000000000110110000100100000000000000000001000100011110101;
ram[ 24 ]= 64'b 0000000000000000110101001101101100000000000000001000111000111001;
ram[ 25 ]= 64'b 0000000000000000110100010100110100000000000000001001001101101000;
ram[ 26 ]= 64'b 0000000000000000110011011001111100000000000000001001100001111111;
ram[ 27 ]= 64'b 0000000000000000110010011101000100000000000000001001110101111111;
ram[ 28 ]= 64'b 0000000000000000110001011110010000000000000000001010001001100111;
ram[ 29 ]= 64'b 0000000000000000110000011101100000000000000000001010011100110110;
ram[ 30 ]= 64'b 0000000000000000101111011010111000000000000000001010101111101011;
ram[ 31 ]= 64'b 0000000000000000101110010110100000000000000000001011000010000101;
ram[ 32 ]= 64'b 0000000000000000101101010000010000000000000000001011010100000100;
ram[ 33 ]= 64'b 0000000000000000101100001000010100000000000000001011100101101000;
ram[ 34 ]= 64'b 0000000000000000101010111110101100000000000000001011110110101110;
ram[ 35 ]= 64'b 0000000000000000101001110011011000000000000000001100000111011000;
ram[ 36 ]= 64'b 0000000000000000101000100110011100000000000000001100010111100100;
ram[ 37 ]= 64'b 0000000000000000100111010111111100000000000000001100100111010001;
ram[ 38 ]= 64'b 0000000000000000100110000111111100000000000000001100110110011111;
ram[ 39 ]= 64'b 0000000000000000100100110110100000000000000000001101000101001101;
ram[ 40 ]= 64'b 0000000000000000100011100011100100000000000000001101010011011011;
ram[ 41 ]= 64'b 0000000000000000100010001111010100000000000000001101100001001000;
ram[ 42 ]= 64'b 0000000000000000100000111001110000000000000000001101101110010100;
ram[ 43 ]= 64'b 0000000000000000011111100010111000000000000000001101111010111110;
ram[ 44 ]= 64'b 0000000000000000011110001010110100000000000000001110000111000101;
ram[ 45 ]= 64'b 0000000000000000011100110001100100000000000000001110010010101010;
ram[ 46 ]= 64'b 0000000000000000011011010111010000000000000000001110011101101011;
ram[ 47 ]= 64'b 0000000000000000011001111011110100000000000000001110101000001001;
ram[ 48 ]= 64'b 0000000000000000011000011111011100000000000000001110110010000011;
ram[ 49 ]= 64'b 0000000000000000010111000010001000000000000000001110111011011000;
ram[ 50 ]= 64'b 0000000000000000010101100011111000000000000000001111000100001001;
ram[ 51 ]= 64'b 0000000000000000010100000100110100000000000000001111001100010100;
ram[ 52 ]= 64'b 0000000000000000010010100101000000000000000000001111010011111010;
ram[ 53 ]= 64'b 0000000000000000010001000100011100000000000000001111011010111010;
ram[ 54 ]= 64'b 0000000000000000001111100011001100000000000000001111100001010011;
ram[ 55 ]= 64'b 0000000000000000001110000001011100000000000000001111100111000111;
ram[ 56 ]= 64'b 0000000000000000001100011111000100000000000000001111101100010100;
ram[ 57 ]= 64'b 0000000000000000001010111100010000000000000000001111110000111011;
ram[ 58 ]= 64'b 0000000000000000001001011001000000000000000000001111110100111010;
ram[ 59 ]= 64'b 0000000000000000000111110101011000000000000000001111111000010011;
ram[ 60 ]= 64'b 0000000000000000000110010001011100000000000000001111111011000100;
ram[ 61 ]= 64'b 0000000000000000000100101101010100000000000000001111111101001110;
ram[ 62 ]= 64'b 0000000000000000000011001000111100000000000000001111111110110001;
ram[ 63 ]= 64'b 0000000000000000000001100100100000000000000000001111111111101100;
ram[ 64 ]= 64'b 0000000000000000000000000000000000000000000000010000000000000000;
ram[ 65 ]= 64'b 1111111111111111111110011011011100000000000000001111111111101100;
ram[ 66 ]= 64'b 1111111111111111111100110111000000000000000000001111111110110001;
ram[ 67 ]= 64'b 1111111111111111111011010010101000000000000000001111111101001110;
ram[ 68 ]= 64'b 1111111111111111111001101110100000000000000000001111111011000100;
ram[ 69 ]= 64'b 1111111111111111111000001010100100000000000000001111111000010011;
ram[ 70 ]= 64'b 1111111111111111110110100110111100000000000000001111110100111010;
ram[ 71 ]= 64'b 1111111111111111110101000011101100000000000000001111110000111011;
ram[ 72 ]= 64'b 1111111111111111110011100000111000000000000000001111101100010100;
ram[ 73 ]= 64'b 1111111111111111110001111110100000000000000000001111100111000111;
ram[ 74 ]= 64'b 1111111111111111110000011100110000000000000000001111100001010011;
ram[ 75 ]= 64'b 1111111111111111101110111011100000000000000000001111011010111010;
ram[ 76 ]= 64'b 1111111111111111101101011010111100000000000000001111010011111010;
ram[ 77 ]= 64'b 1111111111111111101011111011001000000000000000001111001100010100;
ram[ 78 ]= 64'b 1111111111111111101010011100000100000000000000001111000100001001;
ram[ 79 ]= 64'b 1111111111111111101000111101110100000000000000001110111011011000;
ram[ 80 ]= 64'b 1111111111111111100111100000100000000000000000001110110010000011;
ram[ 81 ]= 64'b 1111111111111111100110000100001000000000000000001110101000001001;
ram[ 82 ]= 64'b 1111111111111111100100101000101100000000000000001110011101101011;
ram[ 83 ]= 64'b 1111111111111111100011001110011000000000000000001110010010101010;
ram[ 84 ]= 64'b 1111111111111111100001110101001000000000000000001110000111000101;
ram[ 85 ]= 64'b 1111111111111111100000011101000100000000000000001101111010111110;
ram[ 86 ]= 64'b 1111111111111111011111000110001100000000000000001101101110010100;
ram[ 87 ]= 64'b 1111111111111111011101110000101000000000000000001101100001001000;
ram[ 88 ]= 64'b 1111111111111111011100011100011000000000000000001101010011011011;
ram[ 89 ]= 64'b 1111111111111111011011001001011100000000000000001101000101001101;
ram[ 90 ]= 64'b 1111111111111111011001111000000000000000000000001100110110011111;
ram[ 91 ]= 64'b 1111111111111111011000101000000000000000000000001100100111010001;
ram[ 92 ]= 64'b 1111111111111111010111011001100000000000000000001100010111100100;
ram[ 93 ]= 64'b 1111111111111111010110001100100100000000000000001100000111011000;
ram[ 94 ]= 64'b 1111111111111111010101000001010000000000000000001011110110101110;
ram[ 95 ]= 64'b 1111111111111111010011110111101000000000000000001011100101101000;
ram[ 96 ]= 64'b 1111111111111111010010101111101100000000000000001011010100000100;
ram[ 97 ]= 64'b 1111111111111111010001101001011100000000000000001011000010000101;
ram[ 98 ]= 64'b 1111111111111111010000100101000100000000000000001010101111101011;
ram[ 99 ]= 64'b 1111111111111111001111100010011100000000000000001010011100110110;
ram[ 100 ]= 64'b 1111111111111111001110100001101100000000000000001010001001100111;
ram[ 101 ]= 64'b 1111111111111111001101100010111000000000000000001001110101111111;
ram[ 102 ]= 64'b 1111111111111111001100100110000000000000000000001001100001111111;
ram[ 103 ]= 64'b 1111111111111111001011101011001000000000000000001001001101101000;
ram[ 104 ]= 64'b 1111111111111111001010110010010000000000000000001000111000111001;
ram[ 105 ]= 64'b 1111111111111111001001111011011100000000000000001000100011110101;
ram[ 106 ]= 64'b 1111111111111111001001000110101100000000000000001000001110011100;
ram[ 107 ]= 64'b 1111111111111111001000010100000100000000000000000111111000101110;
ram[ 108 ]= 64'b 1111111111111111000111100011101000000000000000000111100010101101;
ram[ 109 ]= 64'b 1111111111111111000110110101010100000000000000000111001100011001;
ram[ 110 ]= 64'b 1111111111111111000110001001010000000000000000000110110101110100;
ram[ 111 ]= 64'b 1111111111111111000101011111011000000000000000000110011110111101;
ram[ 112 ]= 64'b 1111111111111111000100110111110000000000000000000110000111110111;
ram[ 113 ]= 64'b 1111111111111111000100010010011100000000000000000101110000100010;
ram[ 114 ]= 64'b 1111111111111111000011101111011000000000000000000101011000111110;
ram[ 115 ]= 64'b 1111111111111111000011001110101100000000000000000101000001001101;
ram[ 116 ]= 64'b 1111111111111111000010110000010100000000000000000100101001010000;
ram[ 117 ]= 64'b 1111111111111111000010010100010100000000000000000100010001000111;
ram[ 118 ]= 64'b 1111111111111111000001111010110000000000000000000011111000110011;
ram[ 119 ]= 64'b 1111111111111111000001100011100000000000000000000011100000010111;
ram[ 120 ]= 64'b 1111111111111111000001001110101100000000000000000011000111110001;
ram[ 121 ]= 64'b 1111111111111111000000111100010000000000000000000010101111000100;
ram[ 122 ]= 64'b 1111111111111111000000101100010100000000000000000010010110010000;
ram[ 123 ]= 64'b 1111111111111111000000011110110000000000000000000001111101010110;
ram[ 124 ]= 64'b 1111111111111111000000010011101100000000000000000001100100010111;
ram[ 125 ]= 64'b 1111111111111111000000001011000100000000000000000001001011010101;
ram[ 126 ]= 64'b 1111111111111111000000000100111000000000000000000000110010001111;
ram[ 127 ]= 64'b 1111111111111111000000000001001100000000000000000000011001001000;
ram[ 128 ]= 64'b 1111111111111111000000000000000000000000000000000000000000000000;
ram[ 129 ]= 64'b 1111111111111111000000000001001111111111111111111111100110110111;
ram[ 130 ]= 64'b 1111111111111111000000000100111011111111111111111111001101110000;
ram[ 131 ]= 64'b 1111111111111111000000001011000111111111111111111110110100101010;
ram[ 132 ]= 64'b 1111111111111111000000010011101111111111111111111110011011101000;
ram[ 133 ]= 64'b 1111111111111111000000011110110011111111111111111110000010101001;
ram[ 134 ]= 64'b 1111111111111111000000101100010111111111111111111101101001101111;
ram[ 135 ]= 64'b 1111111111111111000000111100010011111111111111111101010000111011;
ram[ 136 ]= 64'b 1111111111111111000001001110101111111111111111111100111000001110;
ram[ 137 ]= 64'b 1111111111111111000001100011100011111111111111111100011111101000;
ram[ 138 ]= 64'b 1111111111111111000001111010110011111111111111111100000111001100;
ram[ 139 ]= 64'b 1111111111111111000010010100010111111111111111111011101110111000;
ram[ 140 ]= 64'b 1111111111111111000010110000010111111111111111111011010110101111;
ram[ 141 ]= 64'b 1111111111111111000011001110101111111111111111111010111110110010;
ram[ 142 ]= 64'b 1111111111111111000011101111011011111111111111111010100111000001;
ram[ 143 ]= 64'b 1111111111111111000100010010011111111111111111111010001111011101;
ram[ 144 ]= 64'b 1111111111111111000100110111110011111111111111111001111000001000;
ram[ 145 ]= 64'b 1111111111111111000101011111011011111111111111111001100001000010;
ram[ 146 ]= 64'b 1111111111111111000110001001010011111111111111111001001010001011;
ram[ 147 ]= 64'b 1111111111111111000110110101010111111111111111111000110011100110;
ram[ 148 ]= 64'b 1111111111111111000111100011101011111111111111111000011101010010;
ram[ 149 ]= 64'b 1111111111111111001000010100000111111111111111111000000111010001;
ram[ 150 ]= 64'b 1111111111111111001001000110101111111111111111110111110001100011;
ram[ 151 ]= 64'b 1111111111111111001001111011011111111111111111110111011100001010;
ram[ 152 ]= 64'b 1111111111111111001010110010010011111111111111110111000111000110;
ram[ 153 ]= 64'b 1111111111111111001011101011001011111111111111110110110010010111;
ram[ 154 ]= 64'b 1111111111111111001100100110000011111111111111110110011110000000;
ram[ 155 ]= 64'b 1111111111111111001101100010111011111111111111110110001010000000;
ram[ 156 ]= 64'b 1111111111111111001110100001101111111111111111110101110110011000;
ram[ 157 ]= 64'b 1111111111111111001111100010011111111111111111110101100011001001;
ram[ 158 ]= 64'b 1111111111111111010000100101000111111111111111110101010000010100;
ram[ 159 ]= 64'b 1111111111111111010001101001011111111111111111110100111101111010;
ram[ 160 ]= 64'b 1111111111111111010010101111101111111111111111110100101011111011;
ram[ 161 ]= 64'b 1111111111111111010011110111101011111111111111110100011010010111;
ram[ 162 ]= 64'b 1111111111111111010101000001010011111111111111110100001001010001;
ram[ 163 ]= 64'b 1111111111111111010110001100100111111111111111110011111000100111;
ram[ 164 ]= 64'b 1111111111111111010111011001100011111111111111110011101000011011;
ram[ 165 ]= 64'b 1111111111111111011000101000000011111111111111110011011000101110;
ram[ 166 ]= 64'b 1111111111111111011001111000000011111111111111110011001001100000;
ram[ 167 ]= 64'b 1111111111111111011011001001011111111111111111110010111010110010;
ram[ 168 ]= 64'b 1111111111111111011100011100011011111111111111110010101100100100;
ram[ 169 ]= 64'b 1111111111111111011101110000101011111111111111110010011110110111;
ram[ 170 ]= 64'b 1111111111111111011111000110001111111111111111110010010001101011;
ram[ 171 ]= 64'b 1111111111111111100000011101000111111111111111110010000101000001;
ram[ 172 ]= 64'b 1111111111111111100001110101001011111111111111110001111000111010;
ram[ 173 ]= 64'b 1111111111111111100011001110011011111111111111110001101101010101;
ram[ 174 ]= 64'b 1111111111111111100100101000101111111111111111110001100010010100;
ram[ 175 ]= 64'b 1111111111111111100110000100001011111111111111110001010111110110;
ram[ 176 ]= 64'b 1111111111111111100111100000100011111111111111110001001101111100;
ram[ 177 ]= 64'b 1111111111111111101000111101110111111111111111110001000100100111;
ram[ 178 ]= 64'b 1111111111111111101010011100000111111111111111110000111011110110;
ram[ 179 ]= 64'b 1111111111111111101011111011001011111111111111110000110011101011;
ram[ 180 ]= 64'b 1111111111111111101101011010111111111111111111110000101100000101;
ram[ 181 ]= 64'b 1111111111111111101110111011100011111111111111110000100101000101;
ram[ 182 ]= 64'b 1111111111111111110000011100110011111111111111110000011110101100;
ram[ 183 ]= 64'b 1111111111111111110001111110100011111111111111110000011000111000;
ram[ 184 ]= 64'b 1111111111111111110011100000111011111111111111110000010011101011;
ram[ 185 ]= 64'b 1111111111111111110101000011101111111111111111110000001111000100;
ram[ 186 ]= 64'b 1111111111111111110110100110111111111111111111110000001011000101;
ram[ 187 ]= 64'b 1111111111111111111000001010100111111111111111110000000111101100;
ram[ 188 ]= 64'b 1111111111111111111001101110100011111111111111110000000100111011;
ram[ 189 ]= 64'b 1111111111111111111011010010101011111111111111110000000010110001;
ram[ 190 ]= 64'b 1111111111111111111100110111000011111111111111110000000001001110;
ram[ 191 ]= 64'b 1111111111111111111110011011011111111111111111110000000000010011;
ram[ 192 ]= 64'b 1111111111111111111111111111111111111111111111110000000000000000;
ram[ 193 ]= 64'b 0000000000000000000001100100100011111111111111110000000000010011;
ram[ 194 ]= 64'b 0000000000000000000011001000111111111111111111110000000001001110;
ram[ 195 ]= 64'b 0000000000000000000100101101010111111111111111110000000010110001;
ram[ 196 ]= 64'b 0000000000000000000110010001011111111111111111110000000100111011;
ram[ 197 ]= 64'b 0000000000000000000111110101011011111111111111110000000111101100;
ram[ 198 ]= 64'b 0000000000000000001001011001000011111111111111110000001011000101;
ram[ 199 ]= 64'b 0000000000000000001010111100010011111111111111110000001111000100;
ram[ 200 ]= 64'b 0000000000000000001100011111000111111111111111110000010011101011;
ram[ 201 ]= 64'b 0000000000000000001110000001011111111111111111110000011000111000;
ram[ 202 ]= 64'b 0000000000000000001111100011001111111111111111110000011110101100;
ram[ 203 ]= 64'b 0000000000000000010001000100011111111111111111110000100101000101;
ram[ 204 ]= 64'b 0000000000000000010010100101000011111111111111110000101100000101;
ram[ 205 ]= 64'b 0000000000000000010100000100110111111111111111110000110011101011;
ram[ 206 ]= 64'b 0000000000000000010101100011111011111111111111110000111011110110;
ram[ 207 ]= 64'b 0000000000000000010111000010001011111111111111110001000100100111;
ram[ 208 ]= 64'b 0000000000000000011000011111011111111111111111110001001101111100;
ram[ 209 ]= 64'b 0000000000000000011001111011110111111111111111110001010111110110;
ram[ 210 ]= 64'b 0000000000000000011011010111010011111111111111110001100010010100;
ram[ 211 ]= 64'b 0000000000000000011100110001100111111111111111110001101101010101;
ram[ 212 ]= 64'b 0000000000000000011110001010110111111111111111110001111000111010;
ram[ 213 ]= 64'b 0000000000000000011111100010111011111111111111110010000101000001;
ram[ 214 ]= 64'b 0000000000000000100000111001110011111111111111110010010001101011;
ram[ 215 ]= 64'b 0000000000000000100010001111010111111111111111110010011110110111;
ram[ 216 ]= 64'b 0000000000000000100011100011100111111111111111110010101100100100;
ram[ 217 ]= 64'b 0000000000000000100100110110100011111111111111110010111010110010;
ram[ 218 ]= 64'b 0000000000000000100110000111111111111111111111110011001001100000;
ram[ 219 ]= 64'b 0000000000000000100111010111111111111111111111110011011000101110;
ram[ 220 ]= 64'b 0000000000000000101000100110011111111111111111110011101000011011;
ram[ 221 ]= 64'b 0000000000000000101001110011011011111111111111110011111000100111;
ram[ 222 ]= 64'b 0000000000000000101010111110101111111111111111110100001001010001;
ram[ 223 ]= 64'b 0000000000000000101100001000010111111111111111110100011010010111;
ram[ 224 ]= 64'b 0000000000000000101101010000010011111111111111110100101011111011;
ram[ 225 ]= 64'b 0000000000000000101110010110100011111111111111110100111101111010;
ram[ 226 ]= 64'b 0000000000000000101111011010111011111111111111110101010000010100;
ram[ 227 ]= 64'b 0000000000000000110000011101100011111111111111110101100011001001;
ram[ 228 ]= 64'b 0000000000000000110001011110010011111111111111110101110110011000;
ram[ 229 ]= 64'b 0000000000000000110010011101000111111111111111110110001010000000;
ram[ 230 ]= 64'b 0000000000000000110011011001111111111111111111110110011110000000;
ram[ 231 ]= 64'b 0000000000000000110100010100110111111111111111110110110010010111;
ram[ 232 ]= 64'b 0000000000000000110101001101101111111111111111110111000111000110;
ram[ 233 ]= 64'b 0000000000000000110110000100100011111111111111110111011100001010;
ram[ 234 ]= 64'b 0000000000000000110110111001010011111111111111110111110001100011;
ram[ 235 ]= 64'b 0000000000000000110111101011111011111111111111111000000111010001;
ram[ 236 ]= 64'b 0000000000000000111000011100010111111111111111111000011101010010;
ram[ 237 ]= 64'b 0000000000000000111001001010101011111111111111111000110011100110;
ram[ 238 ]= 64'b 0000000000000000111001110110101111111111111111111001001010001011;
ram[ 239 ]= 64'b 0000000000000000111010100000100111111111111111111001100001000010;
ram[ 240 ]= 64'b 0000000000000000111011001000001111111111111111111001111000001000;
ram[ 241 ]= 64'b 0000000000000000111011101101100011111111111111111010001111011101;
ram[ 242 ]= 64'b 0000000000000000111100010000100111111111111111111010100111000001;
ram[ 243 ]= 64'b 0000000000000000111100110001010011111111111111111010111110110010;
ram[ 244 ]= 64'b 0000000000000000111101001111101011111111111111111011010110101111;
ram[ 245 ]= 64'b 0000000000000000111101101011101011111111111111111011101110111000;
ram[ 246 ]= 64'b 0000000000000000111110000101001111111111111111111100000111001100;
ram[ 247 ]= 64'b 0000000000000000111110011100011111111111111111111100011111101000;
ram[ 248 ]= 64'b 0000000000000000111110110001010011111111111111111100111000001110;
ram[ 249 ]= 64'b 0000000000000000111111000011101111111111111111111101010000111011;
ram[ 250 ]= 64'b 0000000000000000111111010011101011111111111111111101101001101111;
ram[ 251 ]= 64'b 0000000000000000111111100001001111111111111111111110000010101001;
ram[ 252 ]= 64'b 0000000000000000111111101100010011111111111111111110011011101000;
ram[ 253 ]= 64'b 0000000000000000111111110100111011111111111111111110110100101010;
ram[ 254 ]= 64'b 0000000000000000111111111011000111111111111111111111001101110000;
ram[ 255 ]= 64'b 0000000000000000111111111110110011111111111111111111100110110111;

end


always @(posedge Clk) 
	begin
	if (En)
		begin
		if (We_A)
			ram[Addr_A] <= DI_A;
		DO_A <= ram[Addr_A];
		end
	if (En)
		begin
		if (We_B)
			ram[Addr_B] <= DI_B;
		DO_B <= ram[Addr_B];
		end 
	end


endmodule


